../../../src/spi_controller.sv