../../../src/sd_controller.sv